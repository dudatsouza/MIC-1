library verilog;
use verilog.vl_types.all;
entity bank_regs_vlg_vec_tst is
end bank_regs_vlg_vec_tst;
