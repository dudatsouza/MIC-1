library verilog;
use verilog.vl_types.all;
entity register_4bit_vlg_vec_tst is
end register_4bit_vlg_vec_tst;
