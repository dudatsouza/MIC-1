library verilog;
use verilog.vl_types.all;
entity Shifter_vlg_vec_tst is
end Shifter_vlg_vec_tst;
